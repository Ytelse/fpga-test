module Bram(
    output[3:0] io_out,
    input [3:0] io_in
);



  assign io_out = io_in;
endmodule

